// This file is intentionally left empty.
// The tt_um_NeuroCore top module is defined in project.v.
// See project.v for the TT wrapper that instantiates neurocore_field_sensor.
